`timescale 1ns / 1ps
`default_nettype none

module half_adder(input wire a,
                input wire b,
                output logic s0, 
                output logic c0);

        assign s0 = a ^ b;
        assign c0 = a & b;
endmodule

module full_adder(input wire a,
                input wire b,
                output logic cin,
                output logic s0,
                output logic c0);

        assign s0 = a ^ b ^ cin;
        assign c0 = (a & b) | (b & cin) | (a & cin);
endmodule

module wallace_tree_128_bit (
        input wire clk_in,
        input wire rst_in,
        input wire [127:0] input_1,
        input wire [127:0] input_2,
        output logic output_ready,
        output logic [255:0] squared_output
        );


        logic [127:0] pp [127:0];

        for (int i = 0; i < 128; i++) begin
                assign pp[i] = (input_2[i] == 1'b1) ? input_1 : 128'b0;
        end

        // stage 1

        logic [250:0] i1; // (128 - 2) * 2 - 1 = 251
        logic [250:0] c1;

        half_adder ha (.a(pp[0][2]), .b(pp[1][1]), .sum(i1[0]), .carry(c1[0]));                         // 3
        full_adder fa (.a(pp[0][3]), .b(pp[1][2]), .cin(pp[2][1]) .sum(i1[1]), .carry(c1[1]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[2]));
        half_adder ha (.a(pp[0][5]), .b(pp[1][4]), .sum(i1[0]), .carry(c1[3]));                         // 5
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[4]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[5]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[6]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[7]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[8]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[9]));
        half_adder ha (.a(pp[0][5]), .b(pp[1][4]), .sum(i1[0]), .carry(c1[10]));                        // 8
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[11]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[12]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[13]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[14]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[15]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[16]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[17]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[18]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[19]));
        half_adder ha (.a(pp[0][5]), .b(pp[1][4]), .sum(i1[0]), .carry(c1[20]));                        // 11
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[21]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[22]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[23]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[24]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[25]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[26]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[27]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[28]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[29]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[30]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[31]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[32]));
        half_adder ha (.a(pp[0][5]), .b(pp[1][4]), .sum(i1[0]), .carry(c1[33]));                        // 14
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[34]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[35]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[36]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[37]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[38]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[39]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[40]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[41]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[42]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[43]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[44]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[45]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[46]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[47]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[48]));
        half_adder ha (.a(pp[0][5]), .b(pp[1][4]), .sum(i1[0]), .carry(c1[49]));                         // 17
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[50]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[51]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[52]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[53]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[54]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[55]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[56]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[57]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[58]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[59]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[60]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[61]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[62]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[63]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[64]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[65]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[66]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[67]));
        half_adder ha (.a(pp[0][5]), .b(pp[1][4]), .sum(i1[0]), .carry(c1[68]));                        // 20
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[69]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[70]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        half_adder ha (.a(pp[0][5]), .b(pp[1][4]), .sum(i1[0]), .carry(c1[0]));                         // 23
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        half_adder ha (.a(pp[0][5]), .b(pp[1][4]), .sum(i1[0]), .carry(c1[0]));                         // 26
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        half_adder ha (.a(pp[0][5]), .b(pp[1][4]), .sum(i1[0]), .carry(c1[0]));                         // 29
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        half_adder ha (.a(pp[0][5]), .b(pp[1][4]), .sum(i1[0]), .carry(c1[0]));                         // 32
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        half_adder ha (.a(pp[0][5]), .b(pp[1][4]), .sum(i1[0]), .carry(c1[0]));                         // 35
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        half_adder ha (.a(pp[0][5]), .b(pp[1][4]), .sum(i1[0]), .carry(c1[0]));                         // 38
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        half_adder ha (.a(pp[0][5]), .b(pp[1][4]), .sum(i1[0]), .carry(c1[0]));                         // 41
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        half_adder ha (.a(pp[0][5]), .b(pp[1][4]), .sum(i1[0]), .carry(c1[0]));                         // 44
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        half_adder ha (.a(pp[0][5]), .b(pp[1][4]), .sum(i1[0]), .carry(c1[0]));                         // 47
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        half_adder ha (.a(pp[0][5]), .b(pp[1][4]), .sum(i1[0]), .carry(c1[0]));                         // 50
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        half_adder ha (.a(pp[0][5]), .b(pp[1][4]), .sum(i1[0]), .carry(c1[0]));                         // 53
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        half_adder ha (.a(pp[0][5]), .b(pp[1][4]), .sum(i1[0]), .carry(c1[0]));                         // 56
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        half_adder ha (.a(pp[0][5]), .b(pp[1][4]), .sum(i1[0]), .carry(c1[0]));                         // 59
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        half_adder ha (.a(pp[0][5]), .b(pp[1][4]), .sum(i1[0]), .carry(c1[0]));                         // 62
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        half_adder ha (.a(pp[0][5]), .b(pp[1][4]), .sum(i1[0]), .carry(c1[0]));                         // 66
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        half_adder ha (.a(pp[0][5]), .b(pp[1][4]), .sum(i1[0]), .carry(c1[0]));                         // 69
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        half_adder ha (.a(pp[0][5]), .b(pp[1][4]), .sum(i1[0]), .carry(c1[0]));                         // 72
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        half_adder ha (.a(pp[0][5]), .b(pp[1][4]), .sum(i1[0]), .carry(c1[0]));                         // 75
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        half_adder ha (.a(pp[0][5]), .b(pp[1][4]), .sum(i1[0]), .carry(c1[0]));                         // 78


        half_adder ha (.a(pp[0][5]), .b(pp[1][4]), .sum(i1[0]), .carry(c1[0]));                         // 120
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        half_adder ha (.a(pp[0][5]), .b(pp[1][4]), .sum(i1[0]), .carry(c1[0]));                         // 123
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));
        full_adder fa (.a(pp[0][4]), .b(pp[1][3]), .cin(pp[2][2]) .sum(i1[0]), .carry(c1[0]));          // 125
        

endmodule

`default_nettype wire